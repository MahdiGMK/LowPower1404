.title "Karatsuba CIRC"

* supply voltages
.global Vss Vdd
Vgnd Vgnd 0 DC 0
Vpwr Vpwr 0 DC 3
* Vss Vss Vpwr DC 0
* Vdd Vdd 0 DC 3
Rgnd Vgnd Vss 0.001
Rpwr Vpwr Vmeasin 0.001
Vmeasin Vmeasin Vdd DC 0

* simple transistor model
.MODEL cmosn NMOS LEVEL=1 VT0=0.7 KP=110U GAMMA=0.4 LAMBDA=0.04 PHI=0.7
.MODEL cmosp PMOS LEVEL=1 VT0=-0.7 KP=50U GAMMA=0.57 LAMBDA=0.05 PHI=0.8

* load design and library
.include yosys/prim_cells_cmos.mod
.include bench.mod

* input signals
Vclk clk 0 PULSE(0 3 1 0.1 0.1 0.8 2)
Vrst rst 0 PULSE(0 3 0.5 0.1 0.1 2.9 40)

Xadder clk rst x0 x1 x2 x3 x4 x5 x6 x7 x8 x9 x10 x11 x12 x13 x14 x15 x16 MCCBench

.tran 0.1 40
.save i(Vmeasin) v(Vmeasin)
* .save v(Vmeasin)
* .probe p(counter)
* .save counter:power
.control
set filetype=ascii
* run
* plot v(clk) v(x0)/4+10 v(x1)/4+11 v(x2)/4+12 v(x3)/4+13 v(x4)/4+14 v(x5)/4+15 v(x6)/4+16 v(x7)/4+17 i(Vmeasin)+20
* save i(Vmeasin)
* plot v(clk) v(rst)+5 v(en)+10 v(out0)+20 v(out1)+25 v(out2)+30 Vmeasin#branch+40
.endc

.end
